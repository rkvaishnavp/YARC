module programcounter(

);

endmodule