`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/02/2023 11:25:51 PM
// Design Name: 
// Module Name: core
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module core(
    
);

hazard_detection hazard_detection();
control control();
forwarding forwarding();
exeunit exeunit();
registers registers();
immmaker immmaker();
insmmeory insmemory();
datamemory datamemory();

endmodule
